MACRO SRAM_1Kx32cm4bw
  SIZE 184.525 BY 171.70 ;
END SRAM_1Kx32cm4bw

MACRO SRAM_2Kx32cm8bw
  SIZE 318.925 BY 169.195 ;
END SRAM_2Kx32cm8bw

MACRO SRAM_6Kx32cm16bw
  SIZE 587.725 BY 237.295 ;
END SRAM_6Kx32cm16bw

MACRO SRAM_8Kx32cm16bw
  SIZE 587.725 BY 305.395 ;
END SRAM_8Kx32cm16bw

MACRO ROM_10240x32
  SIZE 307.955 BY 317.635 ;
END ROM_10240x32

MACRO DPRAM_1Kx32cm4bw
  SIZE 344.94 BY 182.15 ;
END DPRAM_1Kx32cm4bw

MACRO DPRAM_256x32cm4bw
  SIZE 344.94 BY 79.98 ;
END DPRAM_256x32cm4bw

MACRO REGFILE_16x24cm4bw
  SIZE 136.20 BY 29.00 ;
END REGFILE_16x24cm4bw

MACRO REGFILE_256x32cm4bw
  SIZE 169.80 BY 57.80 ;
END REGFILE_256x32cm4bw

MACRO REGFILE_64x21cm4bw
  SIZE 123.60 BY 33.00 ;
END REGFILE_64x21cm4bw

MACRO ascdhd_flash1mb
  SIZE 1460 BY 1938 ;
END ascdhd_flash1mb

